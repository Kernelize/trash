module hello (A1, B1);

    input A1;
    output B1;

    assign B = A;

endmodule
