module cntr_n();
endmodule
