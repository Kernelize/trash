module clock();

endmodule
